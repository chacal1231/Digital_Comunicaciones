//-- Fichero baudgen.vh

// 12MHz External Clock
//`define B115200 104
//`define B57600  208
//`define B38400  313
//`define B19200  625
//`define B9600   1250
//`define B4800   2500
//`define B2400   5000
//`define B1200   10000
//`define B600    20000
//`define B300    40000

// 50MHz External Clock
`define B115200 434
`define B57600  868
`define B38400  1302
`define B19200  2604
`define B9600   5208
`define B4800   10417
`define B2400   20833
`define B1200   41667
`define B600    83333
`define B300    166667

// 100MHz External Clock
//`define B115200 868
//`define B57600  1736
//`define B38400  2604
//`define B19200  5208
//`define B9600   10417
//`define B4800   20833
//`define B2400   41667
//`define B1200   83333
//`define B600    166667
//`define B300    333333